magic
tech sky130A
timestamp 1768332756
<< nwell >>
rect -350 -250 -50 130
<< nmos >>
rect -210 -400 -195 -300
<< pmos >>
rect -210 -200 -195 0
<< ndiff >>
rect -255 -305 -210 -300
rect -255 -395 -245 -305
rect -225 -395 -210 -305
rect -255 -400 -210 -395
rect -195 -305 -150 -300
rect -195 -395 -180 -305
rect -160 -395 -150 -305
rect -195 -400 -150 -395
<< pdiff >>
rect -255 -5 -210 0
rect -255 -195 -245 -5
rect -225 -195 -210 -5
rect -255 -200 -210 -195
rect -195 -5 -150 0
rect -195 -195 -180 -5
rect -160 -195 -150 -5
rect -195 -200 -150 -195
<< ndiffc >>
rect -245 -395 -225 -305
rect -180 -395 -160 -305
<< pdiffc >>
rect -245 -195 -225 -5
rect -180 -195 -160 -5
<< psubdiff >>
rect -250 -455 -155 -445
rect -250 -480 -230 -455
rect -180 -480 -155 -455
rect -250 -490 -155 -480
<< nsubdiff >>
rect -260 105 -155 110
rect -260 85 -225 105
rect -195 85 -155 105
rect -260 70 -155 85
<< psubdiffcont >>
rect -230 -480 -180 -455
<< nsubdiffcont >>
rect -225 85 -195 105
<< poly >>
rect -210 0 -195 50
rect -210 -230 -195 -200
rect -260 -240 -195 -230
rect -260 -260 -250 -240
rect -230 -260 -195 -240
rect -260 -270 -195 -260
rect -110 -240 -75 -230
rect -110 -260 -100 -240
rect -80 -260 -75 -240
rect -110 -270 -75 -260
rect -210 -300 -195 -270
rect -210 -425 -195 -400
<< polycont >>
rect -250 -260 -230 -240
rect -100 -260 -80 -240
<< locali >>
rect -260 105 -155 110
rect -260 85 -225 105
rect -195 85 -155 105
rect -260 70 -155 85
rect -255 -5 -215 70
rect -255 -195 -245 -5
rect -225 -195 -215 -5
rect -255 -200 -215 -195
rect -190 -5 -150 0
rect -190 -195 -180 -5
rect -160 -195 -150 -5
rect -260 -240 -225 -230
rect -260 -260 -250 -240
rect -230 -260 -225 -240
rect -260 -270 -225 -260
rect -255 -305 -215 -300
rect -255 -395 -245 -305
rect -225 -395 -215 -305
rect -255 -445 -215 -395
rect -190 -305 -150 -195
rect -110 -240 -75 -230
rect -110 -260 -100 -240
rect -80 -260 -75 -240
rect -110 -270 -75 -260
rect -190 -395 -180 -305
rect -160 -395 -150 -305
rect -190 -400 -150 -395
rect -255 -455 -155 -445
rect -255 -480 -230 -455
rect -180 -480 -155 -455
rect -255 -490 -155 -480
rect -255 -495 -215 -490
<< viali >>
rect -220 85 -200 105
rect -250 -260 -230 -240
rect -100 -260 -80 -240
rect -220 -480 -195 -455
<< metal1 >>
rect -485 105 40 115
rect -485 85 -220 105
rect -200 85 40 105
rect -485 70 40 85
rect -425 -240 -225 -230
rect -425 -260 -250 -240
rect -230 -260 -225 -240
rect -425 -270 -225 -260
rect -190 -240 30 -230
rect -190 -260 -100 -240
rect -80 -260 30 -240
rect -190 -270 30 -260
rect -475 -455 50 -440
rect -475 -480 -220 -455
rect -195 -480 50 -455
rect -475 -495 50 -480
<< labels >>
rlabel metal1 -20 75 -15 80 1 vdd
rlabel metal1 -20 -475 -15 -470 1 vss
rlabel metal1 -15 -255 -5 -235 1 out
rlabel metal1 -415 -250 -400 -240 1 in
<< end >>
